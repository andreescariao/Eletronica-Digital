module test();
  always #1ns begin
    $display("Hello World");
  end
endmodule
